`timescale 1ns / 1ps
module lcd (
    input clk_50MHz,          // Clock da placa
    input reset_n,            // Reset ativo baixo (global)
    input system_on,          // 1 = sistema ligado, 0 = desligado (controlado pela CPU)
    input display_enable,     // Pulso de 1 ciclo quando atualizar LCD (após instrução)
    input [2:0] opcode_last,  // Opcode 3 bits da última instrução
    input [3:0] reg_number,   // Número do reg (dest ou src para DISPLAY, 0-15)
    input [15:0] reg_value,   // Valor signed 16 bits
    // Pinos LCD DE2-115
    output reg [7:0] LCD_DATA,
    output reg LCD_RS,        // 0=comando, 1=dado
    output reg LCD_EN,
    output LCD_RW = 1'b0,     // Sempre escrita
    output LCD_ON = 1'b1      // Backlight ligado
);

// Parâmetros de delay (50MHz)
localparam 
    DELAY_15MS = 750_000,    // >15ms
    DELAY_4_1MS = 205_000,   // >4.1ms
    DELAY_100US = 5_000,     // >100us
    DELAY_40US = 2_000,      // >40us para comandos
    DELAY_2MS = 100_000,     // >2ms para clear
    DELAY_1US = 50;          // Para pulse EN high

// Estados da FSM
localparam [5:0]
    OFF = 0,
    POWER_ON = 1,
    WAIT_15MS = 2,
    FUNC_SET1 = 3,
    PULSE_EN = 4,
    WAIT_4_1MS = 5,
    FUNC_SET2 = 6,
    WAIT_100US1 = 7,
    FUNC_SET3 = 8,
    WAIT_100US2 = 9,
    FUNC_SET_FINAL = 10,
    WAIT_1MS1 = 11, 
    DISP_OFF = 12,
    WAIT_1MS2 = 13,
    DISP_CLEAR = 14,
    WAIT_2MS = 15,
    ENTRY_MODE = 16,
    WAIT_1MS3 = 17,
    DISP_ON = 18,
    WAIT_1MS4 = 19,
    IDLE = 20,
    SET_ADDR1 = 21, // Linha 1: 0x80
    WAIT_1MS5 = 22,
    WRITE_CHAR1 = 23,
    WAIT_1MS6 = 24,
    SET_ADDR2 = 25, // Linha 2: 0xC0
    WAIT_1MS7 = 26,
    WRITE_CHAR2 = 27,
    WAIT_1MS8 = 28,
    CLEAR_SCREEN = 29;
    WAIT_40US = 30;

reg [5:0] state = OFF;
reg [19:0] delay_cnt = 0;
reg [4:0] char_index = 0; // 0-15 para cada linha
reg [7:0] line1 [0:15]; // Buffer linha 1: Operação
reg [7:0] line2 [0:15]; // Buffer linha 2: Reg bin + valor
reg write_pending = 0;
reg clear_pending = 0;
reg init_mode = 0; // Flag para init vs CLEAR

// Conversão signed/abs - com handling de -32768
wire signed [15:0] signed_value = reg_value;
reg [15:0] abs_value;
reg negative;
always @(*) begin
    negative = (signed_value < 0);
    if (signed_value == 16'sh8000) begin // -32768
        abs_value = 32768;
    end else begin
        abs_value = negative ? -signed_value : signed_value;
    end
end


// Binário 16-bit unsigned para 5 dígitos BCD (double dabble)
reg [19:0] bcd;  // 5 nibbles (20 bits)
integer i;
always @(*) begin
    bcd = 0;
    for (i = 15; i >= 0; i = i - 1) begin
        if (bcd[3:0] >= 5) bcd[3:0] = bcd[3:0] + 3;
        if (bcd[7:4] >= 5) bcd[7:4] = bcd[7:4] + 3;
        if (bcd[11:8] >= 5) bcd[11:8] = bcd[11:8] + 3;
        if (bcd[15:12] >= 5) bcd[15:12] = bcd[15:12] + 3;
        if (bcd[19:16] >= 5) bcd[19:16] = bcd[19:16] + 3;
        bcd = {bcd[18:0], abs_value[i]};
    end
end

// Monta buffers line1 e line2 baseado em opcode
always @(posedge clk_50MHz) begin
    if (display_enable && state == IDLE) begin
        // Preenche line1 e line2 com espaços por default
        for (i = 0; i <= 15; i = i + 1) begin
            line1[i] = 8'h20; // Espaço
            line2[i] = 8'h20;
        end
        case (opcode_last)
            3'b000: begin // LOAD
                line1[0] = "L"; line1[1] = "O"; line1[2] = "A"; line1[3] = "D";
            end
            3'b001: begin // ADD
                line1[0] = "A"; line1[1] = "D"; line1[2] = "D";
            end
            3'b010: begin // ADDI
                line1[0] = "A"; line1[1] = "D"; line1[2] = "D"; line1[3] = "I";
            end
            3'b011: begin // SUB
                line1[0] = "S"; line1[1] = "U"; line1[2] = "B";
            end
            3'b100: begin // SUBI
                line1[0] = "S"; line1[1] = "U"; line1[2] = "B"; line1[3] = "I";
            end
            3'b101: begin // MUL
                line1[0] = "M"; line1[1] = "U"; line1[2] = "L";
            end
            3'b110: begin // CLEAR
                line1[0] = "C"; line1[1] = "L"; line1[2] = "E"; line1[3] = "A"; line1[4] = "R";
                clear_pending = 1;
                write_pending = 1;
            end
            3'b111: begin // DISPLAY -> "DPL" per exemplo PDF
                line1[0] = "D"; line1[1] = "P"; line1[2] = "L";
            end
        endcase
        
        if (opcode_last != 3'b110) begin // Não CLEAR: preenche line2 com reg + valor
            // Reg number binário (4 bits '0'/'1')
            line2[0] = reg_number[3] ? 8'h31 : 8'h30;
            line2[1] = reg_number[2] ? 8'h31 : 8'h30;
            line2[2] = reg_number[1] ? 8'h31 : 8'h30;
            line2[3] = reg_number[0] ? 8'h31 : 8'h30;
            line2[4] = 8'h20; // Espaço
            line2[5] = negative ? 8'h2D : 8'h2B; // - ou +
            // 5 dígitos BCD
            line2[6] = 8'h30 + bcd[19:16];
            line2[7] = 8'h30 + bcd[15:12];
            line2[8] = 8'h30 + bcd[11:8];
            line2[9] = 8'h30 + bcd[7:4];
            line2[10] = 8'h30 + bcd[3:0];
            write_pending = 1;
            clear_pending = 0;
        end
        char_index <= 0;
    end
end

// FSM principal
always @(posedge clk_50MHz or negedge reset_n) begin
    if (!reset_n) begin
        state <= OFF;
        delay_cnt <= 0;
        LCD_EN <= 0;
        LCD_RS <= 0;
        LCD_DATA <= 8'h00;
        char_index <= 0;
        write_pending <= 0;
        clear_pending <= 0;
        init_mode <= 0;
    end else begin
        if (!system_on) begin
            state <= OFF;
            init_mode <= 0;
        end else begin
				case (state)
					OFF: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h08;  // Display off
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					POWER_ON: begin
                        init_mode <= 1; // Ativa flag init
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_15MS) begin
                            delay_cnt <= 0;
                            state <= FUNC_SET1;
                        end
					end
					FUNC_SET1: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h30;
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					WAIT_4_1MS: begin
						 delay_cnt <= delay_cnt + 1;
						 if (delay_cnt == DELAY_4_1MS) begin
							  delay_cnt <= 0;
							  state <= FUNC_SET2;
						 end
					end
					FUNC_SET2: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h30;
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					WAIT_100US1: begin
						 delay_cnt <= delay_cnt + 1;
						 if (delay_cnt == DELAY_100US) begin
							  delay_cnt <= 0;
							  state <= FUNC_SET3;
						 end
					end
					FUNC_SET3: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h30;
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					WAIT_100US2: begin
						 delay_cnt <= delay_cnt + 1;
						 if (delay_cnt == DELAY_100US) begin
							  delay_cnt <= 0;
							  state <= FUNC_SET_FINAL;
						 end
					end
					FUNC_SET_FINAL: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h38;  // 8-bit, 2 lines, 5x8
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					DISP_OFF: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h08;
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					DISP_ON: begin
                        LCD_RS <= 0;
                        LCD_DATA <= 8'h0C;
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                        init_mode <= 0; // Init completa
                    end
					DISP_CLEAR: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h01;
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					WAIT_1MS1: begin
						 delay_cnt <= delay_cnt + 1;
                            if (delay_cnt == DELAY_2MS) begin
                                delay_cnt <= 0;
                                state <= ENTRY_MODE;
                            if (clear_pending || state veio de init) begin  // Ajuste para não re-init após clear
                                state <= IDLE;  
                            end else begin
                                state <= ENTRY_MODE;
                            end
						 end
					end
					WAIT_2MS: begin
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_2MS) begin
                            delay_cnt <= 0;
                            if (clear_pending || !init_mode) begin // Se CLEAR ou não init, vai IDLE
                                state <= IDLE;
                                clear_pending <= 0;
                            end else begin
                                state <= ENTRY_MODE;
                            end
                        end
                    end
					 
					ENTRY_MODE: begin
						 LCD_RS <= 0;
						 LCD_DATA <= 8'h06;  // Increment, no shift
						 LCD_EN <= 1;
						 state <= PULSE_EN;
					end
					IDLE: begin
                        if (write_pending) begin
                            state <= SET_ADDR1;
                            char_index <= 0;
                        end else if (!system_on) begin
                            state <= OFF;
                        end
                    end
					SET_ADDR1: begin
                        LCD_RS <= 0;
                        LCD_DATA <= 8'h80; // Linha 1
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                    end
					
					WAIT_1MS5: begin
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_1MS) begin
                            delay_cnt <= 0;
                            state <= WRITE_CHAR1;
                        end
                    end
                    WRITE_CHAR1: begin
                        LCD_RS <= 1;
                        LCD_DATA <= line1[char_index];
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                    end
                    WAIT_1MS6: begin
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_1MS) begin
                            delay_cnt <= 0;
                            if (char_index == 15) begin
                                char_index <= 0;
                                state <= SET_ADDR2; // Vai para linha 2
                            end else begin
                                char_index <= char_index + 1;
                                state <= WRITE_CHAR1;
                            end
                        end
                    end
                    SET_ADDR2: begin
                        LCD_RS <= 0;
                        LCD_DATA <= 8'hC0; // Início linha 2
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                    end
                    WAIT_1MS7: begin
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_1MS) begin
                            delay_cnt <= 0;
                            state <= WRITE_CHAR2;
                        end
                    end
                    WRITE_CHAR2: begin
                        LCD_RS <= 1;
                        LCD_DATA <= line2[char_index];
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                    end
                    WAIT_1MS8: begin
                        delay_cnt <= delay_cnt + 1;
                        if (delay_cnt == DELAY_1MS) begin
                            delay_cnt <= 0;
                            if (char_index == 15) begin
                                char_index <= 0;
                                write_pending <= 0;
                                if (clear_pending) begin
                                    state <= CLEAR_SCREEN;
                                end else begin
                                    state <= IDLE;
                                end
                            end else begin
                                char_index <= char_index + 1;
                                state <= WRITE_CHAR2;
                            end
                        end
                    end
					CLEAR_SCREEN: begin
                        LCD_RS <= 0;
                        LCD_DATA <= 8'h01;
                        LCD_EN <= 1;
                        state <= PULSE_EN;
                        clear_pending <= 0;
                    end
                    PULSE_EN: begin
                        LCD_EN <= 0;
                        delay_cnt <= 0;
                        state <= next_state_after_pulse;
                    end
			endcase
    end
end
end

// Adicione esta reg para next after pulse
reg [5:0] next_state_after_pulse;
always @(*) begin
    next_state_after_pulse = state; // Default para evitar latches
    case (state)
        // --- Sequência de Inicialização
        OFF:            next_state_after_pulse = WAIT_15MS;    // Espera estabilizar VCC
        FUNC_SET1:      next_state_after_pulse = WAIT_4_1MS;   // Após 1º 0x30
        FUNC_SET2:      next_state_after_pulse = WAIT_100US1;  // Após 2º 0x30
        FUNC_SET3:      next_state_after_pulse = WAIT_100US2;  // Após 3º 0x30
        FUNC_SET_FINAL: next_state_after_pulse = WAIT_100US1;  // Após 0x38 (Function Set)
        DISP_OFF:       next_state_after_pulse = WAIT_100US1;  // Após 0x08
        DISP_CLEAR:     next_state_after_pulse = WAIT_2MS;     // Clear leva > 1.53ms [cite: 45]
        ENTRY_MODE:     next_state_after_pulse = WAIT_100US1;  // Após 0x06
        DISP_ON:        next_state_after_pulse = IDLE;         // Inicialização completa -> IDLE

        // --- Operações de Escrita (IDLE) ---
        SET_ADDR1:      next_state_after_pulse = WAIT_40US;    // Configura endereço Linha 1
        WRITE_CHAR1:    next_state_after_pulse = WAIT_40US;    // Escreve char Linha 1
        SET_ADDR2:      next_state_after_pulse = WAIT_40US;    // Configura endereço Linha 2
        WRITE_CHAR2:    next_state_after_pulse = WAIT_40US;    // Escreve char Linha 2
        
        // --- Comandos Especiais ---
        CLEAR_SCREEN:   next_state_after_pulse = WAIT_2MS;     // Limpa tela durante operação

        default:        next_state_after_pulse = IDLE;
    endcase
end

endmodule